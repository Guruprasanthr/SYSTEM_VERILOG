module str;
  string A="ffac1234";
  initial begin
    $display(" A=%h",A.atohex);
  end
endmodule


Output:  A = ffac1234
