module str;
  string A= "1234guru";
  initial begin
    $display("A=%d",A.atoi());
  end
endmodule

Output:A=   1234
