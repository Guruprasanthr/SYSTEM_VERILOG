module str;
  string A= "GURUPRASANTH";
  initial begin
    $display("A=%d",A.len);
  end
endmodule


Output: A= 12
